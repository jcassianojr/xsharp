#DEFINE LOCALE_SYSTEM_DEFAULT   2048
#DEFINE LOCALE_USER_DEFAULT     1024
#DEFINE LOCALE_IFIRSTDAYOFWEEK  0x0000100C
#DEFINE S_OK                    0x00000000L
#DEFINE SPI_GETWORKAREA         48
#define WM_KEYDOWN              0x0100
#define WM_KEYUP                0x0101
