#define nCONST_MAX_INTEGER_ACCURACY 15 
#define nCONST_MAX_NUMERIC_ACCURACY 18 
#define nCONST_MAX_NUMERIC_NUMBER 999999999999999
#define BUFLEN 80 
#define MAXLEN 12 
#define ID_MONTH1 3001 
#define ID_MONTH2 3002 
#define ID_MONTH3 3003 
#define ID_MONTH4 3004 
#define ID_MONTH5 3005 
#define ID_MONTH6 3006 
#define ID_MONTH7 3007 
#define ID_MONTH8 3008 
#define ID_MONTH9 3009 
#define ID_MONTH10 3010 
#define ID_MONTH11 3011 
#define ID_MONTH12 3012 
#define LOCALE_SYSTEM_DEFAULT 2048
#define LOCALE_USER_DEFAULT 1024
#define FSEL_ALL 0
#define FSEL_END 3
#define FSEL_HOME 2
#define FSEL_TRIM 1
#define FSEL_TRIMEND 4
#define IDM_CalcSLEContextMenu "CalcSLEContextMenu"
#define IDA_CalcSLEContextMenu "CalcSLEContextMenu"
#define IDM_CalcSLEContextMenu_File_ID 22567
#define IDM_CalcSLEContextMenu_File_Calculator_ID 22568
#define IDM_PEDateSleContextMenu "PEDateSleContextMenu"
#define IDA_PEDateSleContextMenu "PEDateSleContextMenu"
#define IDM_PEDateSleContextMenu_File_ID 22579
#define IDM_PEDateSleContextMenu_File_Today_ID 22580
#define IDM_PEDateSleContextMenu_File_Calendar_ID 22581
